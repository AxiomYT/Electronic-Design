DHCP V2.4.1
R2 1 5 330
R4 1 0 330
R3 1 18 330
R1 1 6 330

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
